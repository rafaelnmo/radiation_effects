
* rafaelnevesnmello@gmail.com 10/05/2018
* Implementacao XOR v2

*-------------------------------------------------------
* Parametros e modelos
*-------------------------------------------------------
.include 16nm_HP.pm
.include fontes.cir
.include circuito.cir

Iset gnd xor EXP (0 10u 4ns 10ps 10ps 200ps)
*Iset xor gnd EXP (0 340u 2ns 10ps 10ps 200ps)


*-------------------------------------------------------
* Declaracao do circuito
*-------------------------------------------------------
Xbuff_a a buff_a vdd1 gnd buffer
Xbuff_b b buff_b vdd1 gnd buffer

*Xinv_a buff_a buff_not_a vdd1 gnd inversor
*Xinv_b buff_b buff_not_b vdd1 gnd inversor

Xinv_out xor inv vdd3 gnd buffer

*Xxor_v1 buff_a buff_not_a buff_b buff_not_b xor vdd2 gnd xor_v1
Xxor_v2 buff_a buff_b xor vdd2 gnd xor_v2
*Xxor_v3 buff_a buff_b xor vdd2 gnd xor_v3
*Xxor_v4 buff_a buff_b xor vdd2 gnd xor_v4
*Xxor_v5 buff_a buff_not_a buff_b buff_not_b xor vdd2 gnd xor_v5
*Xxor_v6 buff_a buff_not_a buff_b buff_not_b xor vdd2 gnd xor_v6 
*Xxor_v7 buff_a buff_not_a buff_b buff_not_b xor vdd2 gnd xor_v7
*Xxor_v8 buff_a buff_b xor vdd2 gnd xor_v8
*Xxor_v9 buff_a buff_b buff_not_b xor vdd2 gnd xor_v9
*Xxor_vtest buff_a buff_not_a buff_not_b buff_b xor vdd2 gnd xor_vtest

*-------------------------------------------------------
* Estimulos
*-------------------------------------------------------
.tran 0.01ns 8ns

*-------------------------------------------------------
* Controle
*-------------------------------------------------------
.control
*color0 is background color
*color1 is the grid and the test color
*color 2-15 are for the vectors

*use to output a file with all the mesures
*wrdata "test2" buff_a buff_b xor

set color0=rgb:f/f/f
set color1=rgb:0/0/0
run
.endc

*--------------------------------------------------------
* Fim da declaracao
*--------------------------------------------------------
.end
